LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY CA IS
Port(A,B,C,D,REF,SEL: IN STD_LOGIC_VECTOR (1 DownTo 0);
DISPLAY: OUT STD_LOGIC_VECTOR (6 DownTo 0)
);
END ENTITY;

ARCHITECTURE A_CA OF CA IS
SIGNAL Z: STD_LOGIC_VECTOR (1 DownTo 0);
SIGNAL AUX: STD_LOGIC_VECTOR (2 DownTo 0);
CONSTANT MAYOR: STD_LOGIC_VECTOR (6 DownTo 0):= "0000111";
CONSTANT MENOR: STD_LOGIC_VECTOR (6 DownTo 0):= "0110001";
CONSTANT IGUAL: STD_LOGIC_VECTOR (6 DownTo 0):= "0110111";

BEGIN 
WITH SEL SELECT
Z<= A WHEN "00",
    B WHEN "01",
	C WHEN "10",
	D WHEN OTHERS;

COMP: PROCESS (Z,REF)
BEGIN
IF(Z>REF) THEN 
AUX <= "100";
ELSIF(Z<REF) THEN
AUX <= "010";
ELSE
AUX <= "001";
END IF;
END PROCESS COMP;
DECO: PROCESS (AUX)
BEGIN
CASE AUX IS
WHEN "100" => DISPLAY <= MAYOR;
WHEN "010" => DISPLAY <= MENOR;
WHEN OTHERS => DISPLAY <= IGUAL;
END CASE;
END PROCESS DECO;
END A_CA;